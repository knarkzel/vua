module main

pub fn parse(input string, tokens []string) ? {
	return none
}
