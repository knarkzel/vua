module main

pub fn lex(input string) ? {
	return none
}
