module main

pub fn compile(input string, ast []string) ? {
	return none
}

pub fn eval(program string) ? {
}
